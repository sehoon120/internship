module accumulator (
    input clk, rst, valid_in,
    input [DW-1:0] in_add,
    input [ADDR_WIDTH-1:0] index,  // b*H*P index
    output reg [DW-1:0] y_out,
    output reg valid_out
);



endmodule